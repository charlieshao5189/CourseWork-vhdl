--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   21:26:55 02/04/2016
-- Design Name:   
-- Module Name:   C:/Users/qhsam/Desktop/VHDLv2/smt_watch/dbutton_tb.vhd
-- Project Name:  smt_watch
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: dButton
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY dbutton_tb IS
END dbutton_tb;
 
ARCHITECTURE behavior OF dbutton_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT dButton
    PORT(
         clk : IN  std_logic;
         rst : IN  std_logic;
         btn : IN  std_logic;
         btn_press : OUT  std_logic;
         btn_hold : OUT  std_logic;
         btn_release : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal rst : std_logic := '0';
   signal btn : std_logic := '0';

 	--Outputs
   signal btn_press : std_logic;
   signal btn_hold : std_logic;
   signal btn_release : std_logic;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: dButton PORT MAP (
          clk => clk,
          rst => rst,
          btn => btn,
          btn_press => btn_press,
          btn_hold => btn_hold,
          btn_release => btn_release
        );

  -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   rst_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 800 ns;	
		rst <= '1';
      wait for clk_period;
		rst <= '0';

   end process;
	
   btn_proc: process
   begin		
		wait for clk_period;
		btn <= '1';
		wait for clk_period;
		btn <= not btn;
		wait for clk_period;
		btn <= not btn;
		wait for clk_period;
		btn <= not btn;	
		wait for clk_period;
		btn <= not btn;		
		wait for clk_period;
		btn <= not btn;
		wait for clk_period;
		btn <= not btn;		
      wait for clk_period*12;	
		btn <= not btn;	

   end process;


END;
